library verilog;
use verilog.vl_types.all;
entity AbsSignTestBench is
end AbsSignTestBench;
