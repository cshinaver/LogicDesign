library verilog;
use verilog.vl_types.all;
entity controller is
    generic(
        idle            : integer := 0;
        init            : integer := 1;
        fetch           : integer := 2;
        decode          : integer := 3;
        load            : integer := 4;
        store           : integer := 5;
        add             : integer := 6;
        ldc             : integer := 7;
        sub             : integer := 8;
        jmpz            : integer := 9;
        jmpzjmp         : integer := 10;
        fetch_wait      : integer := 11;
        load_wait       : integer := 12;
        jmp             : integer := 13;
        jmpn            : integer := 14;
        jmpnjmp         : integer := 15;
        loadr           : integer := 16;
        loadr_wait      : integer := 17;
        storer          : integer := 18;
        op_load         : integer := 0;
        op_store        : integer := 1;
        op_add          : integer := 2;
        op_ldc          : integer := 3;
        op_sub          : integer := 4;
        op_jmpz         : integer := 5;
        op_jmp          : integer := 6;
        op_jmpn         : integer := 7;
        op_loadr        : integer := 8;
        op_storer       : integer := 9
    );
    port(
        clk             : in     vl_logic;
        start           : in     vl_logic;
        reset           : in     vl_logic;
        inst            : in     vl_logic_vector(15 downto 0);
        RF_Rp_zero      : in     vl_logic;
        RF_Rp_neg       : in     vl_logic;
        RF_W_addr       : out    vl_logic_vector(3 downto 0);
        RF_W_wr         : out    vl_logic;
        RF_Rp_addr      : out    vl_logic_vector(3 downto 0);
        RF_Rp_rd        : out    vl_logic;
        RF_Rq_addr      : out    vl_logic_vector(3 downto 0);
        RF_Rq_rd        : out    vl_logic;
        PC_clr          : out    vl_logic;
        PC_ld           : out    vl_logic;
        PC_inc          : out    vl_logic;
        I_rd            : out    vl_logic;
        IR_ld           : out    vl_logic;
        D_rd            : out    vl_logic;
        D_wr            : out    vl_logic;
        RF_s1           : out    vl_logic;
        RF_s0           : out    vl_logic;
        alu_s1          : out    vl_logic;
        alu_s0          : out    vl_logic;
        D_addr          : out    vl_logic_vector(7 downto 0);
        RF_W_data       : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of idle : constant is 1;
    attribute mti_svvh_generic_type of init : constant is 1;
    attribute mti_svvh_generic_type of fetch : constant is 1;
    attribute mti_svvh_generic_type of decode : constant is 1;
    attribute mti_svvh_generic_type of load : constant is 1;
    attribute mti_svvh_generic_type of store : constant is 1;
    attribute mti_svvh_generic_type of add : constant is 1;
    attribute mti_svvh_generic_type of ldc : constant is 1;
    attribute mti_svvh_generic_type of sub : constant is 1;
    attribute mti_svvh_generic_type of jmpz : constant is 1;
    attribute mti_svvh_generic_type of jmpzjmp : constant is 1;
    attribute mti_svvh_generic_type of fetch_wait : constant is 1;
    attribute mti_svvh_generic_type of load_wait : constant is 1;
    attribute mti_svvh_generic_type of jmp : constant is 1;
    attribute mti_svvh_generic_type of jmpn : constant is 1;
    attribute mti_svvh_generic_type of jmpnjmp : constant is 1;
    attribute mti_svvh_generic_type of loadr : constant is 1;
    attribute mti_svvh_generic_type of loadr_wait : constant is 1;
    attribute mti_svvh_generic_type of storer : constant is 1;
    attribute mti_svvh_generic_type of op_load : constant is 1;
    attribute mti_svvh_generic_type of op_store : constant is 1;
    attribute mti_svvh_generic_type of op_add : constant is 1;
    attribute mti_svvh_generic_type of op_ldc : constant is 1;
    attribute mti_svvh_generic_type of op_sub : constant is 1;
    attribute mti_svvh_generic_type of op_jmpz : constant is 1;
    attribute mti_svvh_generic_type of op_jmp : constant is 1;
    attribute mti_svvh_generic_type of op_jmpn : constant is 1;
    attribute mti_svvh_generic_type of op_loadr : constant is 1;
    attribute mti_svvh_generic_type of op_storer : constant is 1;
end controller;
