library verilog;
use verilog.vl_types.all;
entity BusMuxTestBench is
end BusMuxTestBench;
